.title KiCad schematic
U7 GND Net-_R13-Pad2_ Net-_R14-Pad1_ Net-_U5-Pad1_ unconnected-_U7-Pad5_ GND unconnected-_U7-Pad7_ +5V NE555P
R13 +5V Net-_R13-Pad2_ R
R14 Net-_R14-Pad1_ Net-_Q1-Pad1_ R
L1 +5V Net-_D3-Pad1_ L
D3 Net-_D3-Pad1_ +5V DIODE
Q1 Net-_Q1-Pad1_ Net-_D3-Pad1_ GND IRLZ34N
R1 Net-_R1-Pad1_ Net-_R1-Pad1_ 10k
R3 Net-_R1-Pad1_ GND 10k
R6 VCC Net-_R6-Pad2_ 10k
R2 Net-_R2-Pad1_ Net-_R2-Pad1_ 10k
R4 Net-_R2-Pad1_ GND 10k
U3 Net-_R5-Pad2_ Net-_R6-Pad2_ Net-_D2-Pad2_ 74HC00
U1 Net-_R5-Pad2_ Net-_R1-Pad1_ unconnected-_U1-Pad3_ LM393
R5 VCC Net-_R5-Pad2_ 10k
U2 Net-_R6-Pad2_ Net-_R2-Pad1_ unconnected-_U2-Pad3_ LM393
U4 Net-_D2-Pad2_ Net-_D1-Pad2_ 74HC04
U6 Net-_R13-Pad2_ Net-_C1-Pad1_ Net-_R11-Pad2_ LM324
C3 Net-_C1-Pad1_ GND 47uF
R9 Net-_D1-Pad2_ Net-_C1-Pad1_ 10k
R11 +5V Net-_R11-Pad2_ 1k
R12 Net-_R11-Pad2_ GND 1k
C1 Net-_C1-Pad1_ GND 47uF
D1 Net-_C1-Pad1_ Net-_D1-Pad2_ DIODE
R7 +5V Net-_R7-Pad2_ 1k
R8 Net-_R7-Pad2_ GND 1k
U5 Net-_U5-Pad1_ Net-_C2-Pad1_ Net-_R7-Pad2_ LM324
R10 Net-_D2-Pad2_ Net-_C2-Pad1_ 20k
D2 Net-_C2-Pad1_ Net-_D2-Pad2_ DIODE
C2 Net-_C2-Pad1_ GND 470uF
.end
